module Decoder_3_to_8 (
    input[0:2] i,
    output[0:7] y
);
and (y[0],i[0],i[1],i[2])

    
endmodule